    Mac OS X            	   2  �     �                                    ATTR;���  �  $  Y                 $   9  com.apple.quarantine   ]     com.apple.lastuseddate#PS E1-  m   5  )com.apple.metadata:kMDItemDownloadedDate   �   �  %com.apple.metadata:kMDItemWhereFroms 0083;5b949c52;Safari;5E02E037-F2C8-43E1-B994-0F1079FE2A19R��[    ��=,    bplist00�3A��i�aq2
                            bplist00�_^https://eee.uci.edu/toolbox/dropbox/download.php/kfarsany_lab2s_tb.vhd?op=getfile&file=5369781_Ihttps://eee.uci.edu/toolbox/dropbox/index.php?op=openfolder&folder=537800l                            �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  This resource fork intentionally left blank                                                                                                                                                                                                                            ��