    Mac OS X            	   2  �     �                                    ATTR;���  �  $  Y                 $   9  com.apple.quarantine   ]     com.apple.lastuseddate#PS 1F-  m   5  )com.apple.metadata:kMDItemDownloadedDate   �   �  %com.apple.metadata:kMDItemWhereFroms 0083;5b949c62;Safari;6A3E680E-F2AE-4C1F-ACDD-CE4B968DF914b��[    :�"    bplist00�3A��i�K��
                            bplist00�_^https://eee.uci.edu/toolbox/dropbox/download.php/kfarsany_lab3s_tb.vhd?op=getfile&file=5371036_Ihttps://eee.uci.edu/toolbox/dropbox/index.php?op=openfolder&folder=537919l                            �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  This resource fork intentionally left blank                                                                                                                                                                                                                            ��