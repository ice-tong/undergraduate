    Mac OS X            	   2  �     �                                    ATTR;���  �  $  V                 $   9  com.apple.quarantine   ]     com.apple.lastuseddate#PS 0F-  m   5  )com.apple.metadata:kMDItemDownloadedDate   �   �  %com.apple.metadata:kMDItemWhereFroms 0083;5b949c4d;Safari;BCAC5946-5785-4D0F-A4B4-5ABE4BAE3A71M��[    ĝ�     bplist00�3A��i�ț�
                            bplist00�_[https://eee.uci.edu/toolbox/dropbox/download.php/kfarsany_lab2b.vhd?op=getfile&file=5369418_Ihttps://eee.uci.edu/toolbox/dropbox/index.php?op=openfolder&folder=537798i                            �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     This resource fork intentionally left blank                                                                                                                                                                                                                            ��