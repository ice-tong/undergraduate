    Mac OS X            	   2  �     �                                    ATTR;���  �  $  V                 $   9  com.apple.quarantine   ]     com.apple.lastuseddate#PS 2F-  m   5  )com.apple.metadata:kMDItemDownloadedDate   �   �  %com.apple.metadata:kMDItemWhereFroms 0083;5b949c3d;Safari;08FB9530-CA53-462F-85F0-898AB55951A3=��[    O
�4    bplist00�3A��i��U�
                            bplist00�_[https://eee.uci.edu/toolbox/dropbox/download.php/kfarsany_lab1s.vhd?op=getfile&file=5368885_Ihttps://eee.uci.edu/toolbox/dropbox/index.php?op=openfolder&folder=537545i                            �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     This resource fork intentionally left blank                                                                                                                                                                                                                            ��