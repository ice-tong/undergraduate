    Mac OS X            	   2  �     �                                    ATTR;���  �  $  V                 $   9  com.apple.quarantine   ]     com.apple.lastuseddate#PS 6E-  m   5  )com.apple.metadata:kMDItemDownloadedDate   �   �  %com.apple.metadata:kMDItemWhereFroms 0083;5b949c6c;Safari;69DFD766-A7F7-4A6E-8AF4-B7C9DF7634B3l��[    �ǝ    bplist00�3A��i�(&�
                            bplist00�_[https://eee.uci.edu/toolbox/dropbox/download.php/kfarsany_lab4s.vhd?op=getfile&file=5374212_Ihttps://eee.uci.edu/toolbox/dropbox/index.php?op=openfolder&folder=538049i                            �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     This resource fork intentionally left blank                                                                                                                                                                                                                            ��