    Mac OS X            	   2  �     �                                    ATTR;���  �  $  V                 $   9  com.apple.quarantine   ]     com.apple.lastuseddate#PS DA-  m   5  )com.apple.metadata:kMDItemDownloadedDate   �   �  %com.apple.metadata:kMDItemWhereFroms 0083;5b949c51;Safari;8CA8A5CB-1443-41DA-9717-9C8E13A7DBAAQ��[    ��9    bplist00�3A��i��6�
                            bplist00�_[https://eee.uci.edu/toolbox/dropbox/download.php/kfarsany_lab2s.vhd?op=getfile&file=5369780_Ihttps://eee.uci.edu/toolbox/dropbox/index.php?op=openfolder&folder=537800i                            �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     This resource fork intentionally left blank                                                                                                                                                                                                                            ��