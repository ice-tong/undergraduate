    Mac OS X            	   2  �     �                                    ATTR;���  �  $  Z                 $   9  com.apple.quarantine   ]     com.apple.lastuseddate#PS 34-  m   5  )com.apple.metadata:kMDItemDownloadedDate   �   �  %com.apple.metadata:kMDItemWhereFroms 0083;5b949c3c;Safari;E922EEC7-D57B-4134-9213-A84BCE3278DD<��[    D#�.    bplist00�3A��i�f�c
                            bplist00�__https://eee.uci.edu/toolbox/dropbox/download.php/kfarsany_lab_1s_tb.vhd?op=getfile&file=5368887_Ihttps://eee.uci.edu/toolbox/dropbox/index.php?op=openfolder&folder=537545m                            �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                 This resource fork intentionally left blank                                                                                                                                                                                                                            ��