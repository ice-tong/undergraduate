    Mac OS X            	   2  �     �                                    ATTR;���  �  $  Y                 $   9  com.apple.quarantine   ]     com.apple.lastuseddate#PS 96-  m   5  )com.apple.metadata:kMDItemDownloadedDate   �   �  %com.apple.metadata:kMDItemWhereFroms 0083;5b949c6c;Safari;5915300E-DA19-4096-8C9F-A4D9BE8FDFFCl��[    .�4    bplist00�3A��i�t@[
                            bplist00�_^https://eee.uci.edu/toolbox/dropbox/download.php/kfarsany_lab4s_tb.vhd?op=getfile&file=5374213_Ihttps://eee.uci.edu/toolbox/dropbox/index.php?op=openfolder&folder=538049l                            �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  This resource fork intentionally left blank                                                                                                                                                                                                                            ��