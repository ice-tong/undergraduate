    Mac OS X            	   2  �     �                                    ATTR;���  �  $  V                 $   9  com.apple.quarantine   ]     com.apple.lastuseddate#PS E3-  m   5  )com.apple.metadata:kMDItemDownloadedDate   �   �  %com.apple.metadata:kMDItemWhereFroms 0083;5b949c38;Safari;B547ABD1-5AA9-42E3-B97A-74501BB865D68��[    �j    bplist00�3A��i�!)
                            bplist00�_[https://eee.uci.edu/toolbox/dropbox/download.php/kfarsany_lab1b.vhd?op=getfile&file=5368303_Ihttps://eee.uci.edu/toolbox/dropbox/index.php?op=openfolder&folder=537541i                            �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     This resource fork intentionally left blank                                                                                                                                                                                                                            ��