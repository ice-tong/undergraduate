    Mac OS X            	   2  �     �                                    ATTR;���  �  $  Y                 $   9  com.apple.quarantine   ]     com.apple.lastuseddate#PS 1A-  m   5  )com.apple.metadata:kMDItemDownloadedDate   �   �  %com.apple.metadata:kMDItemWhereFroms 0083;5b949c67;Safari;C260048D-5E41-411A-8501-3474DE3C8179g��[    ��t    bplist00�3A��i�I�
                            bplist00�_^https://eee.uci.edu/toolbox/dropbox/download.php/kfarsany_lab4b_tb.vhd?op=getfile&file=5372251_Ihttps://eee.uci.edu/toolbox/dropbox/index.php?op=openfolder&folder=538039l                            �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  This resource fork intentionally left blank                                                                                                                                                                                                                            ��