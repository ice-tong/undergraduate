    Mac OS X            	   2  �     �                                    ATTR;���  �  $  V                 $   9  com.apple.quarantine   ]     com.apple.lastuseddate#PS F3-  m   5  )com.apple.metadata:kMDItemDownloadedDate   �   �  %com.apple.metadata:kMDItemWhereFroms 0083;5b949c58;Safari;84335CC2-0CD9-47F3-ACB2-0CB4B476D142X��[    �M�$    bplist00�3A��i�Q2
                            bplist00�_[https://eee.uci.edu/toolbox/dropbox/download.php/kfarsany_lab3b.vhd?op=getfile&file=5370359_Ihttps://eee.uci.edu/toolbox/dropbox/index.php?op=openfolder&folder=537917i                            �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     This resource fork intentionally left blank                                                                                                                                                                                                                            ��