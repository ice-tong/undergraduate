    Mac OS X            	   2  �     �                                    ATTR;���  �  $  V                 $   9  com.apple.quarantine   ]     com.apple.lastuseddate#PS 49-  m   5  )com.apple.metadata:kMDItemDownloadedDate   �   �  %com.apple.metadata:kMDItemWhereFroms 0083;5b949c66;Safari;7122DA1D-F145-4449-A98A-BD80B6F515E1f��[    �Am    bplist00�3A��i�)�'
                            bplist00�_[https://eee.uci.edu/toolbox/dropbox/download.php/kfarsany_lab4b.vhd?op=getfile&file=5372250_Ihttps://eee.uci.edu/toolbox/dropbox/index.php?op=openfolder&folder=538039i                            �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     This resource fork intentionally left blank                                                                                                                                                                                                                            ��