    Mac OS X            	   2  �     �                                    ATTR;���  �  $  Y                 $   9  com.apple.quarantine   ]     com.apple.lastuseddate#PS EA-  m   5  )com.apple.metadata:kMDItemDownloadedDate   �   �  %com.apple.metadata:kMDItemWhereFroms 0083;5b949c59;Safari;6674AA28-97CA-4BEA-B0FB-73362048C72BY��[    8*3    bplist00�3A��i쩛�
                            bplist00�_^https://eee.uci.edu/toolbox/dropbox/download.php/kfarsany_lab3b_tb.vhd?op=getfile&file=5370360_Ihttps://eee.uci.edu/toolbox/dropbox/index.php?op=openfolder&folder=537917l                            �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  This resource fork intentionally left blank                                                                                                                                                                                                                            ��