    Mac OS X            	   2  �     �                                    ATTR;���  �  $  Y                 $   9  com.apple.quarantine   ]     com.apple.lastuseddate#PS 4B-  m   5  )com.apple.metadata:kMDItemDownloadedDate   �   �  %com.apple.metadata:kMDItemWhereFroms 0083;5b949c38;Safari;90D26104-7AD6-464B-B307-780549D7528F8��[    �75    bplist00�3A��i�t��
                            bplist00�_^https://eee.uci.edu/toolbox/dropbox/download.php/kfarsany_lab1b_tb.vhd?op=getfile&file=5368304_Ihttps://eee.uci.edu/toolbox/dropbox/index.php?op=openfolder&folder=537541l                            �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  This resource fork intentionally left blank                                                                                                                                                                                                                            ��