    Mac OS X            	   2  �     �                                    ATTR;���  �  $  Y                 $   9  com.apple.quarantine   ]     com.apple.lastuseddate#PS F6-  m   5  )com.apple.metadata:kMDItemDownloadedDate   �   �  %com.apple.metadata:kMDItemWhereFroms 0083;5b949c4e;Safari;8F51B708-FE0C-46F6-AD03-E1C0CA870847N��[    �}    bplist00�3A��i�)v�
                            bplist00�_^https://eee.uci.edu/toolbox/dropbox/download.php/kfarsany_lab2b_tb.vhd?op=getfile&file=5369419_Ihttps://eee.uci.edu/toolbox/dropbox/index.php?op=openfolder&folder=537798l                            �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  This resource fork intentionally left blank                                                                                                                                                                                                                            ��