    Mac OS X            	   2  �     �                                    ATTR;���  �  $  Y                 $   9  com.apple.quarantine   ]     com.apple.lastuseddate#PS 79-  m   5  )com.apple.metadata:kMDItemDownloadedDate   �   �  %com.apple.metadata:kMDItemWhereFroms 0083;5b949c61;Safari;29BBC858-D13A-4079-A199-BBE82A8BAFF6a��[    vE@.    bplist00�3A��i��J
                            bplist00�_^https://eee.uci.edu/toolbox/dropbox/download.php/kfarsany_lab3s_v2.vhd?op=getfile&file=5371035_Ihttps://eee.uci.edu/toolbox/dropbox/index.php?op=openfolder&folder=537919l                            �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  This resource fork intentionally left blank                                                                                                                                                                                                                            ��